module top(input logic [3:0] a,
    output logic [3:0] b);
endmodule